module top(input        clk, reset,
           output [31:0] WriteData, DataAdr,
           output        MemWrite);

  wire [31:0] PC, Instr, ReadData;

  riscvpipeline rvpipeline(clk, reset, PC, Instr, MemWrite, DataAdr, WriteData, ReadData);
  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);

  always @(posedge clk) begin
      if (MemWrite) begin
        if (DataAdr == 100 && WriteData == 25) begin
          $display("Simulation succeeded");
          $finish;
        end else if (DataAdr != 96) begin
          $display("Simulation failed");
          $finish;
        end
      end
  end
endmodule