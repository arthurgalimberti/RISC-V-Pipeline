module top(
  input wire clk,
  input wire reset,
  output wire [31:0] WriteData,
  output wire [31:0] DataAdr,
  output wire MemWrite
);

  wire [31:0] PC, Instr, ReadData;

  riscvsingle rvsingle(
    clk, reset, PC, Instr, MemWrite, DataAdr,
    WriteData, ReadData
  );

  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
endmodule

module riscvsingle(
  input wire clk, reset,
  output wire [31:0] PC,
  input wire [31:0] Instr,
  output wire MemWrite,
  output wire [31:0] ALUResult, WriteData,
  input wire [31:0] ReadData
);

  wire ALUSrc, RegWrite, Jump, Zero;
  wire [1:0] ResultSrc, ImmSrc;
  wire [2:0] ALUControl;
  wire PCSrc;

  controller c(
    Instr[6:0], Instr[14:12], Instr[30], Zero,
    ResultSrc, MemWrite, PCSrc,
    ALUSrc, RegWrite, Jump,
    ImmSrc, ALUControl
  );

  datapath dp(
    clk, reset, ResultSrc, PCSrc,
    ALUSrc, RegWrite,
    ImmSrc, ALUControl,
    Zero, PC, Instr,
    ALUResult, WriteData, ReadData
  );
endmodule


